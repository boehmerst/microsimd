   // created by generatebits
   parameter IMEMMAUWIDTH = 120
