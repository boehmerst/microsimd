package tta0_params is
  constant fu_PARAM_LSU_addrw_g : integer := 15;
  constant fu_PARAM_LSU_dataw_g : integer := 32;
  constant fu_DATA_LSU_addrw_g : integer := 18;
  constant fu_DATA_LSU_dataw_g : integer := 32;
  constant fu_VLSU_addrw_g : integer := 32;
  constant fu_VLSU_dataw_g : integer := 32;
end tta0_params;
